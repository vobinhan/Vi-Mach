module bt_4_5(input [3:0] X, output [1:0] A, output GS, output EO);
    assign A[0] = 

endmodule