module and_1()
endmodule